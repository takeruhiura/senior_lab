`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/01/2025 08:11:04 PM
// Design Name: 
// Module Name: ov7670_top_uart
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
/*On the PC side, we'll use a Python script over UART to grab a frame and save it as a BMP.

1. High-level architecture

FPGA side

OV7670 camera
  D0..D7  ──► JA[0..7]         (Nexys4 DDR PMOD JA)
  PCLK    ──► JB[0]
  HREF    ──► JB[1]
  VSYNC   ──► JB[2]
  XCLK    ◄── JB[3]            (generated by FPGA)
  SIOC    ◄── JB[4]            (I²C/SCCB SCL)
  SIOD    ◄─► JB[5]            (I²C/SCCB SDA)
  3V3/GND ──► 3.3V / GND pins

FPGA logic:
clk_100mhz → XCLK / I2C / UART / frame readout
cam_pclk   → frame capture → dual-port BRAM → UART → USB-UART → PC


PC side

USB-UART (from Nexys4 DDR) → Python (pyserial + Pillow) → BMP file

2. Top-level Verilog (ov7670_top_uart.v)

This ties everything together:

100 MHz system clock

OV7670 config over SCCB (I²C-like) 
Massachusetts Institute of Technology
+1

Frame capture into dual-port RAM (Xilinx XPM)

UART streaming of one full frame (e.g., 160×120 grayscale*/



// ov7670_top_uart.v
module ov7670_top_uart (
    input  wire clk_100mhz,
    input  wire resetn,

    // OV7670 camera interface
    output wire cam_xclk,
    output wire cam_scl,
    inout  wire cam_sda,
    input  wire cam_pclk,
    input  wire cam_vsync,
    input  wire cam_href,
    input  wire [7:0] cam_data,   // D0..D7

    // UART
    output wire uart_tx
);
    // =========================================================
    // 1) Generate ~24-25 MHz XCLK from 100 MHz
    // =========================================================
    reg [1:0] div_cnt = 2'd0;
    always @(posedge clk_100mhz)
        div_cnt <= div_cnt + 1'b1;

    // 100 MHz / 4 = 25 MHz (close enough for OV7670 XCLK) :contentReference[oaicite:1]{index=1}
    assign cam_xclk = div_cnt[1];

    // =========================================================
    // 2) Configure OV7670 over SCCB (I2C-like)
    // =========================================================
    wire cfg_done;

    ov7670_config u_cfg (
        .clk        (clk_100mhz),
        .resetn     (resetn),
        .scl        (cam_scl),
        .sda        (cam_sda),
        .config_done(cfg_done)
    );

    // =========================================================
    // 3) Capture one grayscale frame into dual-port BRAM
    //    Example: 160x120 = 19200 bytes
    // =========================================================
    localparam IMG_W = 160;
    localparam IMG_H = 120;
    localparam FRAME_SIZE = IMG_W * IMG_H;  // 19200

    wire        cap_we;
    wire [14:0] cap_waddr;
    wire [7:0]  cap_wdata;
    wire        frame_done_cam;   // pulse in cam_pclk domain

    ov7670_capture #(
        .IMG_W(IMG_W),
        .IMG_H(IMG_H)
    ) u_cap (
        .pclk       (cam_pclk),
        .vsync      (cam_vsync),
        .href       (cam_href),
        .d          (cam_data),
        .cfg_done   (cfg_done),

        .we         (cap_we),
        .waddr      (cap_waddr),
        .wdata      (cap_wdata),
        .frame_done (frame_done_cam)
    );

    // =========================================================
    // 4) Dual-port frame buffer (Xilinx XPM)
    //    Port A: write in camera clock domain
    //    Port B: read in 100 MHz domain (for UART)
    // =========================================================

    wire [7:0] fb_rd_data;
    reg        fb_rd_en  = 1'b0;
    reg [14:0] fb_rd_addr = 15'd0;

    // Xilinx true dual-port RAM; Vivado will infer primitives.
    // For real design, include `xpm_memory_tdpram.v` or let Vivado
    // auto-infer from this style.

    xpm_memory_tdpram #(
        .ADDR_WIDTH_A(15),
        .ADDR_WIDTH_B(15),
        .MEMORY_SIZE (FRAME_SIZE*8), // bits
        .MEMORY_PRIMITIVE("auto"),
        .CLOCKING_MODE("independent_clock"),
        .READ_LATENCY_B(1),
        .WRITE_DATA_WIDTH_A(8),
        .READ_DATA_WIDTH_B (8)
    ) u_fb (
        .clka   (cam_pclk),
        .ena    (1'b1),
        .wea    (cap_we),
        .addra  (cap_waddr),
        .dina   (cap_wdata),
        .douta  (),             // unused

        .clkb   (clk_100mhz),
        .enb    (fb_rd_en),
        .web    (1'b0),
        .addrb  (fb_rd_addr),
        .dinb   (8'd0),
        .doutb  (fb_rd_data),

        .injectsbiterra(1'b0),
        .injectdbiterra(1'b0),
        .sbiterrb(),
        .dbiterrb()
    );

    // =========================================================
    // 5) Cross frame_done_cam into clk_100mhz domain
    // =========================================================
    reg [1:0] sync_fd = 2'b00;
    always @(posedge clk_100mhz or negedge resetn) begin
        if (!resetn)
            sync_fd <= 2'b00;
        else
            sync_fd <= {sync_fd[0], frame_done_cam};
    end

    wire frame_done_sys = sync_fd[0] & ~sync_fd[1]; // rising edge detect

    // =========================================================
    // 6) UART + frame readout controller
    // =========================================================
    wire        uart_busy;
    reg  [7:0]  uart_data = 8'd0;
    reg         uart_send = 1'b0;

    uart_tx_module #(
        .CLK_FREQ (100_000_000),
        .BAUD_RATE(115200)
    ) u_uart (
        .clk    (clk_100mhz),
        .resetn (resetn),
        .data_in(uart_data),
        .send   (uart_send),
        .tx     (uart_tx),
        .busy   (uart_busy)
    );

    // State machine: when a frame is done, stream FRAME_SIZE bytes over UART
    localparam S_IDLE  = 2'd0;
    localparam S_START = 2'd1;
    localparam S_SEND  = 2'd2;
    reg [1:0]  state = S_IDLE;
    reg [14:0] pix_cnt = 15'd0;

    always @(posedge clk_100mhz or negedge resetn) begin
        if (!resetn) begin
            state      <= S_IDLE;
            fb_rd_en   <= 1'b0;
            fb_rd_addr <= 15'd0;
            pix_cnt    <= 15'd0;
            uart_send  <= 1'b0;
            uart_data  <= 8'd0;
        end else begin
            uart_send <= 1'b0; // default

            case (state)
                S_IDLE: begin
                    fb_rd_en <= 1'b0;
                    pix_cnt  <= 15'd0;
                    fb_rd_addr <= 15'd0;
                    if (frame_done_sys) begin
                        state <= S_START;
                    end
                end

                S_START: begin
                    // enable RAM read
                    fb_rd_en   <= 1'b1;
                    fb_rd_addr <= 15'd0;
                    state      <= S_SEND;
                end

                S_SEND: begin
                    if (!uart_busy) begin
                        // fb_rd_data is valid from previous cycle due to latency = 1
                        uart_data <= fb_rd_data;
                        uart_send <= 1'b1;

                        // Prepare next address
                        fb_rd_addr <= fb_rd_addr + 1'b1;
                        pix_cnt    <= pix_cnt + 1'b1;

                        if (pix_cnt == FRAME_SIZE-1) begin
                            state    <= S_IDLE;
                            fb_rd_en <= 1'b0;
                        end
                    end
                end

                default: state <= S_IDLE;
            endcase
        end
    end

endmodule

